module CONECTORFLAGS(ALMOST_EMPTYff0, ALMOST_FULLff0, EMPTYff0, FULLff0, 
ALMOST_EMPTYff1, ALMOST_FULLff1, EMPTYff1, FULLff1,
ALMOST_EMPTYff2, ALMOST_FULLff2, EMPTYff2, FULLff2,
ALMOST_EMPTYff3, ALMOST_FULLff3, EMPTYff3, FULLff3,
ALMOST_EMPTY_OUT, ALMOST_FULL_OUT, EMPTY_OUT, FULL_OUT);

	input ALMOST_EMPTYff0, ALMOST_FULLff0, EMPTYff0, FULLff0;
	input ALMOST_EMPTYff1, ALMOST_FULLff1, EMPTYff1, FULLff1;
	input ALMOST_EMPTYff2, ALMOST_FULLff2, EMPTYff2, FULLff2;
	input ALMOST_EMPTYff3, ALMOST_FULLff3, EMPTYff3, FULLff3;
	output reg [3:0] ALMOST_EMPTY_OUT, ALMOST_FULL_OUT, EMPTY_OUT, FULL_OUT;
	
	always @(*) begin
		FULL_OUT[0] <= FULLff0;
		FULL_OUT[1] <= FULLff1;
		FULL_OUT[2] <= FULLff2;
		FULL_OUT[3] <= FULLff3;
		
		ALMOST_FULL_OUT[0] <= ALMOST_FULLff0;
		ALMOST_FULL_OUT[1] <= ALMOST_FULLff1;
		ALMOST_FULL_OUT[2] <= ALMOST_FULLff2;
		ALMOST_FULL_OUT[3] <= ALMOST_FULLff3;
		
		ALMOST_EMPTY_OUT[0] <= ALMOST_EMPTYff0;
		ALMOST_EMPTY_OUT[1] <= ALMOST_EMPTYff1;
		ALMOST_EMPTY_OUT[2] <= ALMOST_EMPTYff2;
		ALMOST_EMPTY_OUT[3] <= ALMOST_EMPTYff3;
		
		EMPTY_OUT[0] <= EMPTYff0;
		EMPTY_OUT[1] <= EMPTYff1;
		EMPTY_OUT[2] <= EMPTYff2;
		EMPTY_OUT[3] <= EMPTYff3;
	end
endmodule
		