`include "TRANSACTIONLAYER.v"
`include "TransactionProb.v"

module testbench;

	wire CLOCK, RESET, PUSHDATOENTRADA, POPffg/*Viene del probador*/, SET_INIT/*Viene del probador*/, POPDATOCF;
	wire [1:0] IDINPUT, SEL, WEIGHT;
	wire [3:0] DATO_IN;
	wire [31:0] TABLE;
	wire [6:0] TL_IN, TH_IN;
	wire IDLE;
	wire [3:0] PAUSE_STB, CONTINUE_STB, ERROR_FULL;
	wire [3:0] DATO_OUTffg;
	
	TransactionProb GeneradorSenales(CLOCK, RESET ,PUSHDATOENTRADA, IDINPUT, DATO_IN, TL_IN, TH_IN, SEL, TABLE, WEIGHT, POPDATOCF,POPffg, SET_INIT, IDLE, PAUSE_STB, CONTINUE_STB, ERROR_FULL);
	TRANSACTIONLAYER conductual(CLOCK, RESET ,PUSHDATOENTRADA, IDINPUT, DATO_IN, TL_IN, TH_IN, SEL, TABLE, WEIGHT, POPDATOCF,POPffg, SET_INIT, IDLE, PAUSE_STB, CONTINUE_STB, ERROR_FULL, DATO_OUTffg);
endmodule