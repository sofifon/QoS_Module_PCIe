`include "RoundRobin.v"
`include "RoundRobin_p.v"

module probadorRoundRobintb();

input wire [1:0] SELECT;
input wire [1:0] W;
input wire [31:0] TAB;
input wire CLK, ENB;
output wire [3:0] OUT;

probadorrr prr(SELECT, CLK, TAB, W, ENB);
RoundRobin rr(SELECT, CLK, TAB, W, ENB, OUT);


initial 
	begin
	$dumpfile("robin.vcd");
	$dumpvars;
	end

endmodule 
